module mul (
    input  [3:0] A, B,
    output [7:0] product
);
    assign product = A * B;

endmodule

